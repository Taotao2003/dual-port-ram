package htax_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    `include "ram_env.sv"
    
	`include "ram_txn.sv"
	`include "ram_seqr.sv"

    `include "ram_agent.sv"
	`include "ram_driver.sv"
	`include "ram_monitor.sv"
	`include "ram_seqs.sv"
    
endpackage